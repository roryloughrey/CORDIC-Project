module cordic;
	
endmodule