module testbench;
	
	cordic cordic();
	
	initial
		begin
		end
	
endmodule